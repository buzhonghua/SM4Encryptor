../../../../rtl/sbox.sv