../../../../include/sm4_encryptor_pkg.svh