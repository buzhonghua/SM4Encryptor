../../../../driver/AXI_SM4_v1_0.sv