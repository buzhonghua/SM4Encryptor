../../../../rtl/lru_recorder.sv