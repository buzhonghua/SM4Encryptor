module sbox_memory(
  input [7:0] i
  ,output logic [7:0] o
);
  always_comb unique case(i)
    0: o = (8)'(214);
    1: o = (8)'(144);
    2: o = (8)'(233);
    3: o = (8)'(254);
    4: o = (8)'(204);
    5: o = (8)'(225);
    6: o = (8)'(61);
    7: o = (8)'(183);
    8: o = (8)'(22);
    9: o = (8)'(182);
    10: o = (8)'(20);
    11: o = (8)'(194);
    12: o = (8)'(40);
    13: o = (8)'(251);
    14: o = (8)'(44);
    15: o = (8)'(5);
    16: o = (8)'(43);
    17: o = (8)'(103);
    18: o = (8)'(154);
    19: o = (8)'(118);
    20: o = (8)'(42);
    21: o = (8)'(190);
    22: o = (8)'(4);
    23: o = (8)'(195);
    24: o = (8)'(170);
    25: o = (8)'(68);
    26: o = (8)'(19);
    27: o = (8)'(38);
    28: o = (8)'(73);
    29: o = (8)'(134);
    30: o = (8)'(6);
    31: o = (8)'(153);
    32: o = (8)'(156);
    33: o = (8)'(66);
    34: o = (8)'(80);
    35: o = (8)'(244);
    36: o = (8)'(145);
    37: o = (8)'(239);
    38: o = (8)'(152);
    39: o = (8)'(122);
    40: o = (8)'(51);
    41: o = (8)'(84);
    42: o = (8)'(11);
    43: o = (8)'(67);
    44: o = (8)'(237);
    45: o = (8)'(207);
    46: o = (8)'(172);
    47: o = (8)'(98);
    48: o = (8)'(228);
    49: o = (8)'(179);
    50: o = (8)'(28);
    51: o = (8)'(169);
    52: o = (8)'(201);
    53: o = (8)'(8);
    54: o = (8)'(232);
    55: o = (8)'(149);
    56: o = (8)'(128);
    57: o = (8)'(223);
    58: o = (8)'(148);
    59: o = (8)'(250);
    60: o = (8)'(117);
    61: o = (8)'(143);
    62: o = (8)'(63);
    63: o = (8)'(166);
    64: o = (8)'(71);
    65: o = (8)'(7);
    66: o = (8)'(167);
    67: o = (8)'(252);
    68: o = (8)'(243);
    69: o = (8)'(115);
    70: o = (8)'(23);
    71: o = (8)'(186);
    72: o = (8)'(131);
    73: o = (8)'(89);
    74: o = (8)'(60);
    75: o = (8)'(25);
    76: o = (8)'(230);
    77: o = (8)'(133);
    78: o = (8)'(79);
    79: o = (8)'(168);
    80: o = (8)'(104);
    81: o = (8)'(107);
    82: o = (8)'(129);
    83: o = (8)'(178);
    84: o = (8)'(113);
    85: o = (8)'(100);
    86: o = (8)'(218);
    87: o = (8)'(139);
    88: o = (8)'(248);
    89: o = (8)'(235);
    90: o = (8)'(15);
    91: o = (8)'(75);
    92: o = (8)'(112);
    93: o = (8)'(86);
    94: o = (8)'(157);
    95: o = (8)'(53);
    96: o = (8)'(30);
    97: o = (8)'(36);
    98: o = (8)'(14);
    99: o = (8)'(94);
    100: o = (8)'(99);
    101: o = (8)'(88);
    102: o = (8)'(209);
    103: o = (8)'(162);
    104: o = (8)'(37);
    105: o = (8)'(34);
    106: o = (8)'(124);
    107: o = (8)'(59);
    108: o = (8)'(1);
    109: o = (8)'(33);
    110: o = (8)'(120);
    111: o = (8)'(135);
    112: o = (8)'(212);
    113: o = (8)'(0);
    114: o = (8)'(70);
    115: o = (8)'(87);
    116: o = (8)'(159);
    117: o = (8)'(211);
    118: o = (8)'(39);
    119: o = (8)'(82);
    120: o = (8)'(76);
    121: o = (8)'(54);
    122: o = (8)'(2);
    123: o = (8)'(231);
    124: o = (8)'(160);
    125: o = (8)'(196);
    126: o = (8)'(200);
    127: o = (8)'(158);
    128: o = (8)'(234);
    129: o = (8)'(191);
    130: o = (8)'(138);
    131: o = (8)'(210);
    132: o = (8)'(64);
    133: o = (8)'(199);
    134: o = (8)'(56);
    135: o = (8)'(181);
    136: o = (8)'(163);
    137: o = (8)'(247);
    138: o = (8)'(242);
    139: o = (8)'(206);
    140: o = (8)'(249);
    141: o = (8)'(97);
    142: o = (8)'(21);
    143: o = (8)'(161);
    144: o = (8)'(224);
    145: o = (8)'(174);
    146: o = (8)'(93);
    147: o = (8)'(164);
    148: o = (8)'(155);
    149: o = (8)'(52);
    150: o = (8)'(26);
    151: o = (8)'(85);
    152: o = (8)'(173);
    153: o = (8)'(147);
    154: o = (8)'(50);
    155: o = (8)'(48);
    156: o = (8)'(245);
    157: o = (8)'(140);
    158: o = (8)'(177);
    159: o = (8)'(227);
    160: o = (8)'(29);
    161: o = (8)'(246);
    162: o = (8)'(226);
    163: o = (8)'(46);
    164: o = (8)'(130);
    165: o = (8)'(102);
    166: o = (8)'(202);
    167: o = (8)'(96);
    168: o = (8)'(192);
    169: o = (8)'(41);
    170: o = (8)'(35);
    171: o = (8)'(171);
    172: o = (8)'(13);
    173: o = (8)'(83);
    174: o = (8)'(78);
    175: o = (8)'(111);
    176: o = (8)'(213);
    177: o = (8)'(219);
    178: o = (8)'(55);
    179: o = (8)'(69);
    180: o = (8)'(222);
    181: o = (8)'(253);
    182: o = (8)'(142);
    183: o = (8)'(47);
    184: o = (8)'(3);
    185: o = (8)'(255);
    186: o = (8)'(106);
    187: o = (8)'(114);
    188: o = (8)'(109);
    189: o = (8)'(108);
    190: o = (8)'(91);
    191: o = (8)'(81);
    192: o = (8)'(141);
    193: o = (8)'(27);
    194: o = (8)'(175);
    195: o = (8)'(146);
    196: o = (8)'(187);
    197: o = (8)'(221);
    198: o = (8)'(188);
    199: o = (8)'(127);
    200: o = (8)'(17);
    201: o = (8)'(217);
    202: o = (8)'(92);
    203: o = (8)'(65);
    204: o = (8)'(31);
    205: o = (8)'(16);
    206: o = (8)'(90);
    207: o = (8)'(216);
    208: o = (8)'(10);
    209: o = (8)'(193);
    210: o = (8)'(49);
    211: o = (8)'(136);
    212: o = (8)'(165);
    213: o = (8)'(205);
    214: o = (8)'(123);
    215: o = (8)'(189);
    216: o = (8)'(45);
    217: o = (8)'(116);
    218: o = (8)'(208);
    219: o = (8)'(18);
    220: o = (8)'(184);
    221: o = (8)'(229);
    222: o = (8)'(180);
    223: o = (8)'(176);
    224: o = (8)'(137);
    225: o = (8)'(105);
    226: o = (8)'(151);
    227: o = (8)'(74);
    228: o = (8)'(12);
    229: o = (8)'(150);
    230: o = (8)'(119);
    231: o = (8)'(126);
    232: o = (8)'(101);
    233: o = (8)'(185);
    234: o = (8)'(241);
    235: o = (8)'(9);
    236: o = (8)'(197);
    237: o = (8)'(110);
    238: o = (8)'(198);
    239: o = (8)'(132);
    240: o = (8)'(24);
    241: o = (8)'(240);
    242: o = (8)'(125);
    243: o = (8)'(236);
    244: o = (8)'(58);
    245: o = (8)'(220);
    246: o = (8)'(77);
    247: o = (8)'(32);
    248: o = (8)'(121);
    249: o = (8)'(238);
    250: o = (8)'(95);
    251: o = (8)'(62);
    252: o = (8)'(215);
    253: o = (8)'(203);
    254: o = (8)'(57);
    255: o = (8)'(72);
    default: o = 'X;
  endcase
endmodule
