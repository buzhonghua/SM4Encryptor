../../../../driver/AXI_SM4_v1_0_S00_AXI.sv