../../../../rtl/roll_shifter.sv