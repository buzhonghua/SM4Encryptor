../../../../rtl/xor_tree.sv