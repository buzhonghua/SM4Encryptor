// -------------------------------------------------------
// -- sm4_encryptor.svh
// -------------------------------------------------------
// This file defines the constant parameter used for sm4 encryptor.
// -------------------------------------------------------

package sm4_encryptor;

    parameter integer word_width_p = 32;

endpackage
