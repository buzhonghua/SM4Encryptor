// -------------------------------------------------------
// -- axi_wrapper.sv
// -------------------------------------------------------
// AXI-lite interface wrapper for sm4_encryptor
// -------------------------------------------------------

module axi_wrapper(

);


endmodule

