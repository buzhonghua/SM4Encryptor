../../../../rtl/sm4_encryptor.sv