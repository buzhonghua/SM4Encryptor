// -------------------------------------------------------
// -- top.sv
// -------------------------------------------------------
// Top design of the accelerators.
// -------------------------------------------------------


module top(
    input cli_i
    ,input reset_i

);


endmodule
