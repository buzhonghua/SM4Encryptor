../../../../rtl/turn_transform.sv