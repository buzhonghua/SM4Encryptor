../../../../rtl/key_cache.sv